module cevero_dvfs
#()(
    input   logic       clk_i,
    input   logic       rst_ni,
    input   logic       error_i,
    output  logic [2:0] set_voltage,
    output  logic [2:0] set_frequency
);


endmodule
